** Profile: "SCHEMATIC1-bias"  [ D:\geoff\Documents\OneDrive - he2b.be\Ecole 2019 - 2020\Q2\Bureau_Etude\1803 - Banc d_essais Moteur\BANC_ESSAI_ELECTRONIQUE\Simulations\Pspice\essaissimupspice-pspicefiles\schematic1\bias.sim ] 

** Creating circuit file "bias.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of D:\SPB_DATA\cdssetup\OrCAD_PSpice\17.2.0\PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
